//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.02 (64-bit)
//Part Number: GW5AST-LV138PG484AC1/I0
//Device: GW5AST-138
//Device Version: B
//Created Time: Fri Jul 25 23:38:47 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [7:0] ad;

wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO(dout[31:0]),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[7:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 32;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h40000301C000020026000004C0000207C8FFFFFF26000001C0000107C8FFFFFF;
defparam prom_inst_0.INIT_RAM_01 = 256'hE0000000E0000000E0000000E0000000C0000002C0000001E000000081060102;
defparam prom_inst_0.INIT_RAM_02 = 256'hC0020007C0020007C0020007C0020007C0020007C0020007C0020007C0020007;
defparam prom_inst_0.INIT_RAM_03 = 256'hC0020007C0020007C0020007C0020007C0020007C0020007C0020007C0020007;
defparam prom_inst_0.INIT_RAM_04 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_05 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_06 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_07 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_08 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_09 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050000;
defparam prom_inst_0.INIT_RAM_0A = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_0B = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_0C = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_0D = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_0E = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_0F = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_10 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_11 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_12 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_13 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_14 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_15 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_16 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_17 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_18 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_19 = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_1A = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_1B = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_1C = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_1D = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_1E = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;
defparam prom_inst_0.INIT_RAM_1F = 256'hC0050007C0050007C0050007C0050007C0050007C0050007C0050007C0050007;

endmodule //Gowin_pROM
